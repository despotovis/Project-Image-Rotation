`ifndef BRAM_SEQ_1_SV
`define BRAM_SEQ_1_SV

class bram_seq_1 extends bram_base_seq;

    logic [15:0] mask0 = 16'b0000000000000000;
    logic [15:0] mask1 = 16'b0010000000000000;
    logic [15:0] mask2 = 16'b0100000000000000;
    
    logic [7:0] data1[3600] = {8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01010101,
8'b00110101,
8'b00111000,
8'b00111000,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00111000,
8'b00111000,
8'b00110101,
8'b01010101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01001010,
8'b01100001,
8'b01101011,
8'b01101011,
8'b01100001,
8'b01001010,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111111,
8'b01000101,
8'b01000010,
8'b00111101,
8'b01011010,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01011011,
8'b00111101,
8'b01000010,
8'b01000101,
8'b00111111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110111,
8'b00110111,
8'b01000010,
8'b01100011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100011,
8'b01000011,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110110,
8'b00110111,
8'b01000110,
8'b01101100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101101,
8'b01000110,
8'b00110111,
8'b00110111,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111011,
8'b01101000,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101000,
8'b00111011,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110110,
8'b00110111,
8'b00111011,
8'b01001110,
8'b01100011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101001,
8'b01010011,
8'b01000010,
8'b00111011,
8'b01000100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100100,
8'b01001111,
8'b00111011,
8'b00110111,
8'b00110110,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111100,
8'b00110111,
8'b00110111,
8'b01001001,
8'b01101010,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100001,
8'b00111011,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01000100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101011,
8'b01001001,
8'b00110111,
8'b00110111,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01000100,
8'b01101101,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100100,
8'b00111000,
8'b00110111,
8'b01000110,
8'b01100000,
8'b01101011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101101,
8'b01000101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00110111,
8'b01100100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000010,
8'b00110111,
8'b01001110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000011,
8'b00111011,
8'b01000110,
8'b01100010,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100100,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00111111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000100,
8'b01000011,
8'b01101101,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000100,
8'b00110111,
8'b00110111,
8'b00111000,
8'b01011111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00111111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b01000110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101010,
8'b01001111,
8'b00110111,
8'b00111110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000101,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01000110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01001111,
8'b01001111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000110,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00110111,
8'b01011100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01001111,
8'b01000110,
8'b01010001,
8'b01101001,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01011100,
8'b00110111,
8'b00110110,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01001011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000011,
8'b00111011,
8'b01000001,
8'b01010011,
8'b01101001,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00111101,
8'b00110111,
8'b00110111,
8'b00111101,
8'b01100100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01001011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01100010,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111011,
8'b01100000,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101010,
8'b01011111,
8'b01000101,
8'b00110111,
8'b01000001,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01101100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101011,
8'b01100000,
8'b01000110,
8'b00110111,
8'b00111000,
8'b01100100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101101,
8'b01000100,
8'b01000101,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101011,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01101011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101101,
8'b01001101,
8'b00110111,
8'b01000011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101011,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01100010,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101101,
8'b01000111,
8'b01001011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101001,
8'b01010011,
8'b01000010,
8'b00111011,
8'b01000100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01001011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100001,
8'b00111011,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01000100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01001010,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00110111,
8'b01011100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100100,
8'b00111000,
8'b00110111,
8'b01000110,
8'b01100000,
8'b01101011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01011101,
8'b00110111,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01000110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000010,
8'b00110111,
8'b01001101,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01000110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000011,
8'b00111011,
8'b01000110,
8'b01100010,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101100,
8'b01010001,
8'b00111101,
8'b00111100,
8'b01010000,
8'b01101100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000001,
8'b01000011,
8'b01101101,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000101,
8'b00110111,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b00111111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01000100,
8'b00110111,
8'b00110111,
8'b00111000,
8'b01011111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01010000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01010000,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101101,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00111110,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00110111,
8'b01100011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101010,
8'b01001111,
8'b00110111,
8'b00111110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00111100,
8'b00110111,
8'b01001101,
8'b01001100,
8'b00110111,
8'b00111100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100011,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01000101,
8'b01101101,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01001111,
8'b01001111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101100,
8'b01000100,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111100,
8'b00110110,
8'b00110111,
8'b01001000,
8'b01101010,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101011,
8'b01001000,
8'b00110111,
8'b00110110,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110110,
8'b00110111,
8'b00111011,
8'b01001110,
8'b01100100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100011,
8'b01001111,
8'b00111010,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111011,
8'b01101000,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101000,
8'b00111011,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00111010,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01000110,
8'b01101100,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101100,
8'b01000101,
8'b00110111,
8'b00110110,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01000010,
8'b01100011,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01101110,
8'b01100011,
8'b01000010,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00111111,
8'b01000101,
8'b01000001,
8'b00111100,
8'b01011010,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b01011010,
8'b00111101,
8'b01000010,
8'b01000101,
8'b00111110,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110101,
8'b00110100,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110110,
8'b00110100,
8'b00110101,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01010011,
8'b01010011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b01100011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01110100,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01011111,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01110100,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01010010,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00101110,
8'b00111001,
8'b01001101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01000101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b00111001,
8'b01110011,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110100,
8'b00111001,
8'b00110111,
8'b00101111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01101000,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01101000,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01011011,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01011011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01001110,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01001110,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01000001,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01000001,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00110111,
8'b01110001,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110001,
8'b00111000,
8'b00110110,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01100100,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01100100,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01010111,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01010111,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01000011,
8'b01110001,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110101,
8'b01110001,
8'b01000011,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000};

    logic [7:0] data2[3600] = {8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01010101,
8'b00110101,
8'b00111000,
8'b00111000,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00111000,
8'b00111000,
8'b00110101,
8'b01010101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111000,
8'b01101011,
8'b10101001,
8'b11000101,
8'b11000101,
8'b10101000,
8'b01101011,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01001100,
8'b01011110,
8'b01010101,
8'b01000110,
8'b10010111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10010111,
8'b01000110,
8'b01010101,
8'b01011110,
8'b01001100,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110111,
8'b00110111,
8'b01010101,
8'b10101111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10101111,
8'b01010110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110110,
8'b00110111,
8'b01011111,
8'b11000111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001000,
8'b01100000,
8'b00110111,
8'b00110111,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01000001,
8'b10111100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10111100,
8'b01000001,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110110,
8'b00110111,
8'b01000001,
8'b01110111,
8'b10110000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000000,
8'b10000100,
8'b01010011,
8'b01000001,
8'b01011010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10110001,
8'b01111000,
8'b01000010,
8'b00110111,
8'b00110110,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111100,
8'b00110111,
8'b00110111,
8'b01100111,
8'b11000010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10101000,
8'b01000011,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01011011,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000011,
8'b01100111,
8'b00110111,
8'b00110111,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01011011,
8'b11001001,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10110000,
8'b00111011,
8'b00110111,
8'b01011111,
8'b10100101,
8'b11000100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001001,
8'b01011100,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00110111,
8'b10110000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01010011,
8'b00110111,
8'b01110100,
8'b11001011,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011000,
8'b01000001,
8'b01100001,
8'b10101100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10110000,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b01001101,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011011,
8'b01011001,
8'b11001000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011010,
8'b00110111,
8'b00110111,
8'b00111011,
8'b10100010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01001100,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b01100000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000001,
8'b01111001,
8'b00110111,
8'b01001000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011110,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01011111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001011,
8'b01111001,
8'b01111000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00111000,
8'b10011101,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01110110,
8'b01011111,
8'b01111110,
8'b10111111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10011101,
8'b00111000,
8'b00110110,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01101101,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011000,
8'b01000001,
8'b01010011,
8'b10000100,
8'b11000000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01000111,
8'b00110111,
8'b00110111,
8'b01000110,
8'b10110011,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01101100,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b10101010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011010,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01000100,
8'b10100111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000001,
8'b10100011,
8'b01011110,
8'b00110111,
8'b01010011,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10101000,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b11000110,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000100,
8'b10100101,
8'b01011111,
8'b00110111,
8'b00111011,
8'b10110001,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001000,
8'b01011011,
8'b01011100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b11000101,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001010,
8'b01110011,
8'b00110111,
8'b01010111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000100,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b10101010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001000,
8'b01100100,
8'b01101101,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000000,
8'b10000100,
8'b01010011,
8'b01000001,
8'b01011010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10101000,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01101101,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10101000,
8'b01000011,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01011011,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01101010,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00111000,
8'b10011101,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10110000,
8'b00111011,
8'b00110111,
8'b01100000,
8'b10100101,
8'b11000100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10011100,
8'b00111000,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01011111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01010011,
8'b00110111,
8'b01110100,
8'b11001011,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011110,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01100000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011000,
8'b01000001,
8'b01100001,
8'b10101100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001000,
8'b01111100,
8'b01000110,
8'b01000110,
8'b01111100,
8'b11001000,
8'b11001100,
8'b11001100,
8'b11001011,
8'b01010001,
8'b01010110,
8'b11001000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011110,
8'b00110111,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01001101,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01011010,
8'b00110111,
8'b00110111,
8'b00111011,
8'b10100010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01111100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01111100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001011,
8'b11001010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01001011,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00110111,
8'b10110000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000001,
8'b01111001,
8'b00110111,
8'b01001000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b01000110,
8'b00110111,
8'b01011000,
8'b01010111,
8'b00110111,
8'b01000110,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10101110,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01011100,
8'b11001001,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001011,
8'b01111001,
8'b01111000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001000,
8'b01011010,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111100,
8'b00110110,
8'b00110111,
8'b01100101,
8'b11000010,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000010,
8'b01100100,
8'b00110111,
8'b00110110,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110110,
8'b00110111,
8'b01000001,
8'b01110111,
8'b10110000,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10110000,
8'b01110110,
8'b01000000,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01000001,
8'b10111100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10111100,
8'b01000000,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00111010,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01011111,
8'b11000111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11000111,
8'b01011110,
8'b00110111,
8'b00110110,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01010110,
8'b10101110,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b11001100,
8'b10101110,
8'b01010101,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110110,
8'b00110111,
8'b00110111,
8'b01001011,
8'b01011110,
8'b01010011,
8'b01000101,
8'b10010110,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b10010110,
8'b01000110,
8'b01010100,
8'b01011110,
8'b01001011,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110101,
8'b00110100,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110110,
8'b00110100,
8'b00110101,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01100001,
8'b01100001,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b10001000,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b01111011,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b10011111,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b01100101,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00101110,
8'b00111010,
8'b01011101,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b01001110,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b00111010,
8'b10011101,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10011110,
8'b00111011,
8'b00110111,
8'b00101111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b10001010,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10001010,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01110100,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b01110100,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01011101,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b01011110,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01000111,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b01000111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00111000,
8'b10011001,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10011001,
8'b00111000,
8'b00110110,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b10000011,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10000011,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01101101,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b01101101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01001011,
8'b10011001,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10100000,
8'b10011001,
8'b01001011,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000};

    logic [7:0] data3[3600] = {8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01010101,
8'b00110101,
8'b00111000,
8'b00111000,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00111000,
8'b00111000,
8'b00110101,
8'b01010101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01010110,
8'b01111010,
8'b10001011,
8'b10001011,
8'b01111010,
8'b01010110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01000011,
8'b01001110,
8'b01001001,
8'b01000000,
8'b01110000,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01110000,
8'b01000000,
8'b01001001,
8'b01001110,
8'b01000011,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110111,
8'b00110111,
8'b01001001,
8'b01111110,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111110,
8'b01001010,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110110,
8'b00110111,
8'b01001111,
8'b10001100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001101,
8'b01001111,
8'b00110111,
8'b00110111,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111101,
8'b10000110,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10000110,
8'b00111101,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110110,
8'b00110111,
8'b00111101,
8'b01011101,
8'b01111110,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001000,
8'b01100101,
8'b01001000,
8'b00111101,
8'b01001100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111111,
8'b01011101,
8'b00111110,
8'b00110111,
8'b00110110,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111100,
8'b00110111,
8'b00110111,
8'b01010011,
8'b10001001,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111010,
8'b00111110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01001100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001010,
8'b01010011,
8'b00110111,
8'b00110111,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01001100,
8'b10001101,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111111,
8'b00111001,
8'b00110111,
8'b01001111,
8'b01111000,
8'b10001010,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001101,
8'b01001101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00110111,
8'b01111111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001000,
8'b00110111,
8'b01011011,
8'b10001110,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001011,
8'b00111101,
8'b01010000,
8'b01111100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111111,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b01000100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001100,
8'b01001011,
8'b10001101,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001100,
8'b00110111,
8'b00110111,
8'b00111001,
8'b01110111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01000011,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b01001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001000,
8'b01011110,
8'b00110111,
8'b01000001,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001110,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001110,
8'b01011110,
8'b01011101,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00110111,
8'b01110011,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01011101,
8'b01001111,
8'b01100001,
8'b10000111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01110011,
8'b00110111,
8'b00110110,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01010111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001011,
8'b00111101,
8'b01000111,
8'b01100101,
8'b10001000,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01000001,
8'b00110111,
8'b00110111,
8'b01000000,
8'b10000000,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01010110,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01111011,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001100,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111110,
8'b01111001,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001000,
8'b01110111,
8'b01001110,
8'b00110111,
8'b01000111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111010,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10001011,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001010,
8'b01111000,
8'b01001111,
8'b00110111,
8'b00111001,
8'b01111111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001101,
8'b01001100,
8'b01001101,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001011,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10001011,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001110,
8'b01011011,
8'b00110111,
8'b01001010,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001010,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01111011,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001101,
8'b01010001,
8'b01010111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001000,
8'b01100101,
8'b01001000,
8'b00111101,
8'b01001100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111010,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01010111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111010,
8'b00111110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01001100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01010101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00110111,
8'b01110011,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111111,
8'b00111001,
8'b00110111,
8'b01001111,
8'b01111000,
8'b10001010,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01110011,
8'b00110111,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001000,
8'b00110111,
8'b01011011,
8'b10001110,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001110,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001011,
8'b00111101,
8'b01010000,
8'b01111100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001101,
8'b01100000,
8'b01000000,
8'b01000000,
8'b01100000,
8'b10001101,
8'b10001111,
8'b10001111,
8'b10001110,
8'b01000111,
8'b01001010,
8'b10001101,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001110,
8'b00110111,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01000100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01001100,
8'b00110111,
8'b00110111,
8'b00111001,
8'b01110111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01100000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01100000,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001110,
8'b10001110,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01000011,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00110111,
8'b01111110,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001000,
8'b01011110,
8'b00110111,
8'b01000001,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01000000,
8'b00110111,
8'b01111110,
8'b01111101,
8'b00110111,
8'b01000000,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111101,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01001101,
8'b10001101,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001110,
8'b01011110,
8'b01011101,
8'b10001111,
8'b10001111,
8'b10001111,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001101,
8'b01001100,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111100,
8'b00110110,
8'b00110111,
8'b01010010,
8'b10001001,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001001,
8'b01010010,
8'b00110111,
8'b00110110,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110110,
8'b00110111,
8'b00111101,
8'b01011101,
8'b01111111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111110,
8'b01011101,
8'b00111100,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111101,
8'b10000110,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10000110,
8'b00111101,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00111010,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01001111,
8'b10001100,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001100,
8'b01001110,
8'b00110111,
8'b00110110,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b01001001,
8'b01111101,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b10001111,
8'b01111101,
8'b01001001,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110110,
8'b00110111,
8'b00110111,
8'b01000011,
8'b01001110,
8'b01000111,
8'b00111111,
8'b01101111,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b01101111,
8'b01000000,
8'b01001000,
8'b01001110,
8'b01000011,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110101,
8'b00110101,
8'b00110100,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110110,
8'b00110100,
8'b00110101,
8'b00110101,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110100,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10010010,
8'b10010010,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b11100101,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b10111001,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b10001110,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00101110,
8'b00111101,
8'b01111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b01100100,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b00111101,
8'b11111010,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111011,
8'b00111110,
8'b00110111,
8'b00101111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b11010110,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11010110,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10101011,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b10101011,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10000000,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b10000001,
8'b00110111,
8'b00110111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b01010110,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b01010110,
8'b00110111,
8'b00111000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110011,
8'b00110110,
8'b00111000,
8'b11110010,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11110010,
8'b00111001,
8'b00110110,
8'b00110011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b11001000,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11001000,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110111,
8'b00110111,
8'b10011101,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b10011101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00110110,
8'b00110111,
8'b01011101,
8'b11110010,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11111111,
8'b11110010,
8'b01011101,
8'b00110111,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111000,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00111111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00111001,
8'b00110110,
8'b00110110,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110111,
8'b00110110,
8'b00110111,
8'b00110100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000};
   
    int num_of_addrs = 3600; 
   
    `uvm_object_utils (bram_seq_1)
    
    function new(string name = "bram_seq_1");
        super.new(name);
    endfunction
      
    virtual task body();
        `uvm_info(get_type_name(), $sformatf("A bram is being used, %d ", mask0), UVM_NONE)
        
        for(int i = 0; i < num_of_addrs; i++)begin
            //`uvm_info(get_type_name(), $sformatf("Writing to A bram, to addr %d", i), UVM_NONE)
            `uvm_do_with(req, {req.wr == 1; req.data == data1[i]; req.addr == 16'(mask0 | i);});
        end
        
        `uvm_info(get_type_name(), $sformatf("B bram is being used, %d ", mask1), UVM_NONE)
        
        for(int j = 0; j < num_of_addrs; j++)begin
            //`uvm_info(get_type_name(), $sformatf("Writing to A bram, to addr %d", j), UVM_NONE)
            `uvm_do_with(req, {req.wr == 1; req.data == data2[j]; req.addr == 16'(mask1 | j);});
        end
        
        `uvm_info(get_type_name(), $sformatf("C bram is being used, %d ", mask2), UVM_NONE)
        
        for(int k = 0; k < num_of_addrs; k++)begin
            //`uvm_info(get_type_name(), $sformatf("Writing to A bram, to addr %d", k), UVM_NONE)
            `uvm_do_with(req, {req.wr == 1; req.data == data3[k]; req.addr == 16'(mask2 | k);});
        end
        
        //`uvm_do_with(req, {req.wr == 0; req.data == 0; req.addr == 0;});
        
    endtask : body 

endclass : bram_seq_1

`endif