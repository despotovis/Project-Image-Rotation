`include "axil_base_seq.sv"
`include "bram_base_seq.sv"
`include "axil_seq_1.sv"
`include "bram_seq_1.sv"
`include "axil_seq_2.sv"
`include "bram_seq_2.sv"