`include "test_base.sv"
`include "test_simple.sv"