----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/08/2023 03:31:35 PM
-- Design Name: 
-- Module Name: better_ip_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_textio.all;
use STD.textio.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity better_ip_tb is
generic (
        PIXEL_WIDTH : integer := 8;
        FIXED_POINT_WIDTH : positive := 16;
        WIDTH : positive := 8
    );
end better_ip_tb;

architecture Behavioral of better_ip_tb is
signal clk_i : std_logic;
signal rst_i : std_logic;
signal bram_read_enable_s : std_logic;
signal bram_write_enable_s : std_logic;
signal ready_o : STD_LOGIC;
--signal end_o : std_logic;
signal start_i : STD_LOGIC;
signal snoop_io : STD_LOGIC_VECTOR (FIXED_POINT_WIDTH - 1 downto 0);
signal x_s : STD_LOGIC_VECTOR (WIDTH - 1 downto 0);
signal y_s : STD_LOGIC_VECTOR (WIDTH - 1 downto 0);
signal cx_i : STD_LOGIC_VECTOR (WIDTH - 1 downto 0);
signal cy_i : STD_LOGIC_VECTOR (WIDTH - 1 downto 0);
signal sinc_i : STD_LOGIC_VECTOR (FIXED_POINT_WIDTH - 1 downto 0);
signal cosc_i : STD_LOGIC_VECTOR (FIXED_POINT_WIDTH - 1 downto 0);
signal midx_i : STD_LOGIC_VECTOR (WIDTH - 1 downto 0);
signal midy_i : STD_LOGIC_VECTOR (WIDTH - 1 downto 0);
--signal row_i : STD_LOGIC_VECTOR (WIDTH - 1 downto 0);
--signal col_i : STD_LOGIC_VECTOR (WIDTH - 1 downto 0);
signal lr_i  : STD_LOGIC;
 signal new_heigth_i :  STD_LOGIC_VECTOR(WIDTH - 1 downto 0 );
  signal new_width_i :  STD_LOGIC_VECTOR(WIDTH - 1 downto 0 );
  signal old_width_i :  STD_LOGIC_VECTOR(WIDTH - 1 downto 0 ); 
  signal old_heigth_i :  STD_LOGIC_VECTOR(WIDTH - 1 downto 0 );
  signal row_s :  STD_LOGIC_VECTOR(WIDTH - 1 downto 0 );
  signal col_s :   STD_LOGIC_VECTOR(WIDTH - 1 downto 0 );
 --signal x_i:  STD_LOGIC_VECTOR(WIDTH - 1 downto 0 );
 -- signal y_i :   STD_LOGIC_VECTOR(WIDTH - 1 downto 0 );
  signal calc_req_s:  STD_LOGIC; 
  signal calc_finished_s :  STD_LOGIC;
  signal calc_ready_s : STD_LOGIC;
  signal pixel_data_r_in :  STD_LOGIC_VECTOR(PIXEL_WIDTH - 1 downto 0);
  signal pixel_data_g_in :  STD_LOGIC_VECTOR(PIXEL_WIDTH - 1 downto 0);
  signal pixel_data_b_in :  STD_LOGIC_VECTOR(PIXEL_WIDTH - 1 downto 0);
  signal pixel_address_unrotated1_o :  STD_LOGIC_VECTOR (2*WIDTH - 1 downto 0);
  signal pixel_data_r_o :  STD_LOGIC_VECTOR(PIXEL_WIDTH - 1 downto 0);
  signal pixel_data_g_o :  STD_LOGIC_VECTOR(PIXEL_WIDTH - 1 downto 0);
  signal pixel_data_b_o :  STD_LOGIC_VECTOR(PIXEL_WIDTH - 1 downto 0);
  signal pixel_address_rotated1_o :  STD_LOGIC_VECTOR (2*WIDTH - 1 downto 0);
  
  type inputDataT is array (0 to 3599) of std_logic_vector(7 downto 0);
  type outputDataT is array (0 to 7055) of std_logic_vector(7 downto 0);
  
  --shared variable fstatus : file_open_status;
  --file output1 : text;
  shared variable L : line;
  
  file output1 : text is out "C:\Users\micac\Desktop\PSDS project\o_r.txt";
  --file output2 : text; --is out "C:\Users\micac\Desktop\PSDS project\o_g.txt";
  --file output3 : text; --is out "C:\Users\micac\Desktop\PSDS project\o_b.txt";
  
  shared variable inputDataR : inputDataT := 
  (
  "00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01010101",
"00110101",
"00111000",
"00111000",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00111000",
"00111000",
"00110101",
"01010101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110111",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"01001010",
"01100001",
"01101011",
"01101011",
"01100001",
"01001010",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"00110111",
"00111111",
"01000101",
"01000010",
"00111101",
"01011010",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01011011",
"00111101",
"01000010",
"01000101",
"00111111",
"00110111",
"00110111",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110111",
"00110111",
"01000010",
"01100011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100011",
"01000011",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110110",
"00110111",
"01000110",
"01101100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101101",
"01000110",
"00110111",
"00110111",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"00111011",
"01101000",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101000",
"00111011",
"00110111",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110110",
"00110111",
"00111011",
"01001110",
"01100011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101001",
"01010011",
"01000010",
"00111011",
"01000100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100100",
"01001111",
"00111011",
"00110111",
"00110110",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110111",
"00110111",
"01001001",
"01101010",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100001",
"00111011",
"00110111",
"00110111",
"00110111",
"01000100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101011",
"01001001",
"00110111",
"00110111",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01000100",
"01101101",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100100",
"00111000",
"00110111",
"01000110",
"01100000",
"01101011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101101",
"01000101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00110111",
"01100100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000010",
"00110111",
"01001110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000011",
"00111011",
"01000110",
"01100010",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100100",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00111111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000100",
"01000011",
"01101101",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000100",
"00110111",
"00110111",
"00111000",
"01011111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"00111111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"01000110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101010",
"01001111",
"00110111",
"00111110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000101",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01000110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01001111",
"01001111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000110",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00110111",
"01011100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01001111",
"01000110",
"01010001",
"01101001",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01011100",
"00110111",
"00110110",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01001011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000011",
"00111011",
"01000001",
"01010011",
"01101001",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"00111101",
"00110111",
"00110111",
"00111101",
"01100100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01001011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01100010",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000100",
"00110111",
"00110111",
"00110111",
"00111011",
"01100000",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101010",
"01011111",
"01000101",
"00110111",
"01000001",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100001",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01101100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101011",
"01100000",
"01000110",
"00110111",
"00111000",
"01100100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101101",
"01000100",
"01000101",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101011",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01101011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101101",
"01001101",
"00110111",
"01000011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101011",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01100010",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101101",
"01000111",
"01001011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101001",
"01010011",
"01000010",
"00111011",
"01000100",
"01101110",
"01101110",
"01101110",
"01101110",
"01100001",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01001011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100001",
"00111011",
"00110111",
"00110111",
"00110111",
"01000100",
"01101110",
"01101110",
"01101110",
"01101110",
"01001010",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00110111",
"01011100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100100",
"00111000",
"00110111",
"01000110",
"01100000",
"01101011",
"01101110",
"01101110",
"01101110",
"01101110",
"01011101",
"00110111",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01000110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000010",
"00110111",
"01001101",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01000110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000011",
"00111011",
"01000110",
"01100010",
"01101110",
"01101110",
"01101110",
"01101110",
"01101100",
"01010001",
"00111101",
"00111100",
"01010000",
"01101100",
"01101110",
"01101110",
"01101110",
"01000001",
"01000011",
"01101101",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000101",
"00110111",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"00111111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01000100",
"00110111",
"00110111",
"00111000",
"01011111",
"01101110",
"01101110",
"01101110",
"01010000",
"00110111",
"00110111",
"00110111",
"00110111",
"01010000",
"01101110",
"01101110",
"01101110",
"01101110",
"01101101",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"00111110",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00110111",
"01100011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101010",
"01001111",
"00110111",
"00111110",
"01101110",
"01101110",
"01101110",
"00111100",
"00110111",
"01001101",
"01001100",
"00110111",
"00111100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100011",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01000101",
"01101101",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01001111",
"01001111",
"01101110",
"01101110",
"01101110",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101100",
"01000100",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110110",
"00110111",
"01001000",
"01101010",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101011",
"01001000",
"00110111",
"00110110",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110110",
"00110111",
"00111011",
"01001110",
"01100100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100011",
"01001111",
"00111010",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"00111011",
"01101000",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101000",
"00111011",
"00110111",
"00110111",
"00110110",
"00111010",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"01000110",
"01101100",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01101100",
"01000101",
"00110111",
"00110110",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"01000010",
"01100011",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"01101110",
"01101110",
"01101110",
"01101110",
"01101110",
"01100011",
"01000010",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110110",
"00110111",
"00110111",
"00111111",
"01000101",
"01000001",
"00111100",
"01011010",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"01011010",
"00111101",
"01000010",
"01000101",
"00111110",
"00110111",
"00110111",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110111",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110101",
"00110100",
"00110110",
"00110110",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"00110110",
"00110110",
"00110100",
"00110101",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01010011",
"01010011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"01100011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01110100",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01011111",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01110100",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01010010",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00101110",
"00111001",
"01001101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01000101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"00111001",
"01110011",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110100",
"00111001",
"00110111",
"00101111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01101000",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01101000",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01011011",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01011011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01001110",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01001110",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01000001",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01000001",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00110111",
"01110001",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110001",
"00111000",
"00110110",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01100100",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01100100",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01010111",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01010111",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01000011",
"01110001",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110101",
"01110001",
"01000011",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
  ); 
  
  shared variable inputDataG : inputDataT :=
  (
  "00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01010101",
"00110101",
"00111000",
"00111000",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00111000",
"00111000",
"00110101",
"01010101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110111",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00111000",
"01101011",
"10101001",
"11000101",
"11000101",
"10101000",
"01101011",
"00111000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"00110111",
"01001100",
"01011110",
"01010101",
"01000110",
"10010111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10010111",
"01000110",
"01010101",
"01011110",
"01001100",
"00110111",
"00110111",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110111",
"00110111",
"01010101",
"10101111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10101111",
"01010110",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110110",
"00110111",
"01011111",
"11000111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001000",
"01100000",
"00110111",
"00110111",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"01000001",
"10111100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10111100",
"01000001",
"00110111",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110110",
"00110111",
"01000001",
"01110111",
"10110000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000000",
"10000100",
"01010011",
"01000001",
"01011010",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10110001",
"01111000",
"01000010",
"00110111",
"00110110",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110111",
"00110111",
"01100111",
"11000010",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10101000",
"01000011",
"00110111",
"00110111",
"00110111",
"01011011",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000011",
"01100111",
"00110111",
"00110111",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01011011",
"11001001",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10110000",
"00111011",
"00110111",
"01011111",
"10100101",
"11000100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001001",
"01011100",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00110111",
"10110000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01010011",
"00110111",
"01110100",
"11001011",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011000",
"01000001",
"01100001",
"10101100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10110000",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"01001101",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011011",
"01011001",
"11001000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011010",
"00110111",
"00110111",
"00111011",
"10100010",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01001100",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"01100000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000001",
"01111001",
"00110111",
"01001000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011110",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01011111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001011",
"01111001",
"01111000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00111000",
"10011101",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01110110",
"01011111",
"01111110",
"10111111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10011101",
"00111000",
"00110110",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01101101",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011000",
"01000001",
"01010011",
"10000100",
"11000000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01000111",
"00110111",
"00110111",
"01000110",
"10110011",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01101100",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"10101010",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011010",
"00110111",
"00110111",
"00110111",
"01000100",
"10100111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000001",
"10100011",
"01011110",
"00110111",
"01010011",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10101000",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"11000110",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000100",
"10100101",
"01011111",
"00110111",
"00111011",
"10110001",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001000",
"01011011",
"01011100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"11000101",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001010",
"01110011",
"00110111",
"01010111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000100",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"10101010",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001000",
"01100100",
"01101101",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000000",
"10000100",
"01010011",
"01000001",
"01011010",
"11001100",
"11001100",
"11001100",
"11001100",
"10101000",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01101101",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10101000",
"01000011",
"00110111",
"00110111",
"00110111",
"01011011",
"11001100",
"11001100",
"11001100",
"11001100",
"01101010",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00111000",
"10011101",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10110000",
"00111011",
"00110111",
"01100000",
"10100101",
"11000100",
"11001100",
"11001100",
"11001100",
"11001100",
"10011100",
"00111000",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01011111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01010011",
"00110111",
"01110100",
"11001011",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011110",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01100000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011000",
"01000001",
"01100001",
"10101100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001000",
"01111100",
"01000110",
"01000110",
"01111100",
"11001000",
"11001100",
"11001100",
"11001011",
"01010001",
"01010110",
"11001000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011110",
"00110111",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01001101",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01011010",
"00110111",
"00110111",
"00111011",
"10100010",
"11001100",
"11001100",
"11001100",
"01111100",
"00110111",
"00110111",
"00110111",
"00110111",
"01111100",
"11001100",
"11001100",
"11001100",
"11001011",
"11001010",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"01001011",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00110111",
"10110000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000001",
"01111001",
"00110111",
"01001000",
"11001100",
"11001100",
"11001100",
"01000110",
"00110111",
"01011000",
"01010111",
"00110111",
"01000110",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10101110",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01011100",
"11001001",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001011",
"01111001",
"01111000",
"11001100",
"11001100",
"11001100",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001000",
"01011010",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110110",
"00110111",
"01100101",
"11000010",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000010",
"01100100",
"00110111",
"00110110",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110110",
"00110111",
"01000001",
"01110111",
"10110000",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10110000",
"01110110",
"01000000",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"01000001",
"10111100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10111100",
"01000000",
"00110111",
"00110111",
"00110110",
"00111010",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"01011111",
"11000111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"11000111",
"01011110",
"00110111",
"00110110",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"01010110",
"10101110",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"11001100",
"11001100",
"11001100",
"11001100",
"11001100",
"10101110",
"01010101",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110110",
"00110111",
"00110111",
"01001011",
"01011110",
"01010011",
"01000101",
"10010110",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"10010110",
"01000110",
"01010100",
"01011110",
"01001011",
"00110111",
"00110111",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110111",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"00111000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110101",
"00110100",
"00110110",
"00110110",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"00110110",
"00110110",
"00110100",
"00110101",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01100001",
"01100001",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"10001000",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"01111011",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"10011111",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"01100101",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00101110",
"00111010",
"01011101",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"01001110",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"00111010",
"10011101",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10011110",
"00111011",
"00110111",
"00101111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"10001010",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10001010",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01110100",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"01110100",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01011101",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"01011110",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01000111",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"01000111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00111000",
"10011001",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10011001",
"00111000",
"00110110",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"10000011",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10000011",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01101101",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"01101101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01001011",
"10011001",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10100000",
"10011001",
"01001011",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
  );
  
  shared variable inputDataB : inputDataT :=
  (
  "00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01010101",
"00110101",
"00111000",
"00111000",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00111000",
"00111000",
"00110101",
"01010101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110111",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"01010110",
"01111010",
"10001011",
"10001011",
"01111010",
"01010110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"00110111",
"01000011",
"01001110",
"01001001",
"01000000",
"01110000",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01110000",
"01000000",
"01001001",
"01001110",
"01000011",
"00110111",
"00110111",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110111",
"00110111",
"01001001",
"01111110",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111110",
"01001010",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110110",
"00110111",
"01001111",
"10001100",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001101",
"01001111",
"00110111",
"00110111",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"00111101",
"10000110",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10000110",
"00111101",
"00110111",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110110",
"00110111",
"00111101",
"01011101",
"01111110",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001000",
"01100101",
"01001000",
"00111101",
"01001100",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111111",
"01011101",
"00111110",
"00110111",
"00110110",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110111",
"00110111",
"01010011",
"10001001",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111010",
"00111110",
"00110111",
"00110111",
"00110111",
"01001100",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001010",
"01010011",
"00110111",
"00110111",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01001100",
"10001101",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111111",
"00111001",
"00110111",
"01001111",
"01111000",
"10001010",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001101",
"01001101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00110111",
"01111111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001000",
"00110111",
"01011011",
"10001110",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001011",
"00111101",
"01010000",
"01111100",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111111",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"01000100",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001100",
"01001011",
"10001101",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001100",
"00110111",
"00110111",
"00111001",
"01110111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01000011",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"01001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001000",
"01011110",
"00110111",
"01000001",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001110",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001110",
"01011110",
"01011101",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00110111",
"01110011",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01011101",
"01001111",
"01100001",
"10000111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01110011",
"00110111",
"00110110",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01010111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001011",
"00111101",
"01000111",
"01100101",
"10001000",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01000001",
"00110111",
"00110111",
"01000000",
"10000000",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01010110",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01111011",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001100",
"00110111",
"00110111",
"00110111",
"00111110",
"01111001",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001000",
"01110111",
"01001110",
"00110111",
"01000111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111010",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10001011",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001010",
"01111000",
"01001111",
"00110111",
"00111001",
"01111111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001101",
"01001100",
"01001101",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001011",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10001011",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001110",
"01011011",
"00110111",
"01001010",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001010",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01111011",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001101",
"01010001",
"01010111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001000",
"01100101",
"01001000",
"00111101",
"01001100",
"10001111",
"10001111",
"10001111",
"10001111",
"01111010",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01010111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111010",
"00111110",
"00110111",
"00110111",
"00110111",
"01001100",
"10001111",
"10001111",
"10001111",
"10001111",
"01010101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00110111",
"01110011",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111111",
"00111001",
"00110111",
"01001111",
"01111000",
"10001010",
"10001111",
"10001111",
"10001111",
"10001111",
"01110011",
"00110111",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001000",
"00110111",
"01011011",
"10001110",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001110",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001011",
"00111101",
"01010000",
"01111100",
"10001111",
"10001111",
"10001111",
"10001111",
"10001101",
"01100000",
"01000000",
"01000000",
"01100000",
"10001101",
"10001111",
"10001111",
"10001110",
"01000111",
"01001010",
"10001101",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001110",
"00110111",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01000100",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01001100",
"00110111",
"00110111",
"00111001",
"01110111",
"10001111",
"10001111",
"10001111",
"01100000",
"00110111",
"00110111",
"00110111",
"00110111",
"01100000",
"10001111",
"10001111",
"10001111",
"10001110",
"10001110",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01000011",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00110111",
"01111110",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001000",
"01011110",
"00110111",
"01000001",
"10001111",
"10001111",
"10001111",
"01000000",
"00110111",
"01111110",
"01111101",
"00110111",
"01000000",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111101",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01001101",
"10001101",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001110",
"01011110",
"01011101",
"10001111",
"10001111",
"10001111",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001101",
"01001100",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111100",
"00110110",
"00110111",
"01010010",
"10001001",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001001",
"01010010",
"00110111",
"00110110",
"00111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110110",
"00110111",
"00111101",
"01011101",
"01111111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111110",
"01011101",
"00111100",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"00111101",
"10000110",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10000110",
"00111101",
"00110111",
"00110111",
"00110110",
"00111010",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"01001111",
"10001100",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001100",
"01001110",
"00110111",
"00110110",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"01001001",
"01111101",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"10001111",
"10001111",
"10001111",
"10001111",
"10001111",
"01111101",
"01001001",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110110",
"00110111",
"00110111",
"01000011",
"01001110",
"01000111",
"00111111",
"01101111",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"01101111",
"01000000",
"01001000",
"01001110",
"01000011",
"00110111",
"00110111",
"00110110",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110111",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110101",
"00110101",
"00110100",
"00110110",
"00110110",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"00110110",
"00110110",
"00110100",
"00110101",
"00110101",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110100",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10010010",
"10010010",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"11100101",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"10111001",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"10001110",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00101110",
"00111101",
"01111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01100100",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"00111101",
"11111010",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111011",
"00111110",
"00110111",
"00101111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"11010110",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11010110",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10101011",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"10101011",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10000000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"10000001",
"00110111",
"00110111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"01010110",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"01010110",
"00110111",
"00111000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110011",
"00110110",
"00111000",
"11110010",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11110010",
"00111001",
"00110110",
"00110011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"11001000",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11001000",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110111",
"00110111",
"10011101",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"10011101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00110110",
"00110111",
"01011101",
"11110010",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11111111",
"11110010",
"01011101",
"00110111",
"00110110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111000",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00111001",
"00110110",
"00110110",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110111",
"00110110",
"00110111",
"00110100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
  );
  
  shared variable outputDataR : outputDataT := (others => (others => '0'));
  shared variable outputDataG : outputDataT := (others => (others => '0'));
  shared variable outputDataB : outputDataT := (others => (others => '0'));
  
begin
fsm: entity work.rot_fsm
    generic map (PIXEL_WIDTH => PIXEL_WIDTH,
                 FIXED_POINT_WIDTH => FIXED_POINT_WIDTH,
                 WIDTH => WIDTH)
    port map (clk_i => clk_i,
              rst_i => rst_i,
              bram_read_enable_o => bram_read_enable_s,
              bram_write_enable_o => bram_write_enable_s,
              ready_o => ready_o,
              --end_o => end_o,
              start_i => start_i,
              new_heigth_i => new_heigth_i,
              new_width_i => new_width_i,
              old_width_i => old_width_i,
              old_heigth_i => old_heigth_i,
              row_o => row_s,
              col_o => col_s,
              x_i => x_s,
              y_i => y_s,
              calc_req_o => calc_req_s,
              calc_finished_i => calc_finished_s,
              calc_ready_i => calc_ready_s,
              pixel_data_r_in => pixel_data_r_in,
              pixel_data_g_in =>  pixel_data_g_in,
              pixel_data_b_in =>  pixel_data_b_in,
              pixel_address_unrotated1_o => pixel_address_unrotated1_o,
              pixel_data_r_o => pixel_data_r_o,
              pixel_data_g_o =>  pixel_data_g_o,
              pixel_data_b_o =>  pixel_data_b_o,
              pixel_address_rotated1_o => pixel_address_rotated1_o
              );
pru: entity work.point_rotation_unit 
    generic map (FIXED_POINT_WIDTH => FIXED_POINT_WIDTH,
                 WIDTH => WIDTH)
    port map (clk_i => clk_i,
              rst_i => rst_i,
              ready_o => calc_ready_s,
              start => calc_req_s,
              finished_o => calc_finished_S,
              snoop_io => snoop_io,
              x_o => x_s,
              y_o => y_s,
              cx_i => cx_i,
              cy_i => cy_i,
              sinc_i => sinc_i,
              cosc_i => cosc_i,
              midx_i => midx_i,
              midy_i => midy_i,
              row_i => row_s,
              col_i => col_s,
              lr_i =>  lr_i
              );
              
    pixelDataR : process(bram_read_enable_s, pixel_address_unrotated1_o)
    begin
        if(bram_read_enable_s = '1') then
            pixel_data_r_in <= inputDataR(TO_INTEGER(unsigned(pixel_address_unrotated1_o)));
        end if;
    end process;
    
    pixelDataG : process(bram_read_enable_s, pixel_address_unrotated1_o)
    begin
        if(bram_read_enable_s = '1') then
            pixel_data_g_in <= inputDataG(TO_INTEGER(unsigned(pixel_address_unrotated1_o)));
        end if;
    end process;
    
    pixelDataB : process(bram_read_enable_s, pixel_address_unrotated1_o)
    begin
        if(bram_read_enable_s = '1') then
            pixel_data_b_in <= inputDataB(TO_INTEGER(unsigned(pixel_address_unrotated1_o)));
        end if;
    end process;
    
    writeDataR : process(bram_write_enable_s, pixel_address_rotated1_o)
    begin
        --file_open(fstatus, output1, "C:\Users\micac\Desktop\PSDS project\o_r.txt", WRITE_MODE);
        if(bram_write_enable_s = '1') then
            outputDataR(TO_INTEGER(unsigned(pixel_address_rotated1_o))) := pixel_data_r_o;
            write(L, pixel_address_rotated1_o);
            writeline(output1, L);
        end if;
    end process;
    
    writeDataG : process(bram_write_enable_s, pixel_address_rotated1_o)
    begin
        if(bram_write_enable_s = '1') then
            outputDataG(TO_INTEGER(unsigned(pixel_address_rotated1_o))) := pixel_data_g_o;
        end if;
    end process;
    
    writeDataB : process(bram_write_enable_s, pixel_address_rotated1_o)
    begin
        if(bram_write_enable_s = '1') then
            outputDataB(TO_INTEGER(unsigned(pixel_address_rotated1_o))) := pixel_data_b_o;
        end if;
    end process;
              
clk: 
    process begin
        clk_i <= '1';
        wait for 50ns;
        clk_i <= '0';
        wait for 50ns;
    end process;
init: process begin
        rst_i <= '1';
        wait for 100ns;
        rst_i <= '0';
        if ready_o /= '1' then
            wait until ready_o = '1';
        end if;
        wait for 100ns; 
        lr_i <= '0';
        new_heigth_i <=std_logic_vector(to_signed(integer( real(84)),WIDTH));
        new_width_i <= std_logic_vector(to_signed(integer( real(84)),WIDTH));
        old_heigth_i <=std_logic_vector(to_signed(integer( real(60)),WIDTH));
        old_width_i <= std_logic_vector(to_signed(integer( real(60)),WIDTH));
        sinc_i <= std_logic_vector(to_signed(integer( real(0.70710678118)*real(2**WIDTH)),FIXED_POINT_WIDTH));
        cosc_i <= std_logic_vector(to_signed(integer( real(0.70710678118)*real(2**WIDTH)),FIXED_POINT_WIDTH));
        cx_i <= std_logic_vector(to_signed(integer( real(30)),WIDTH));
        cy_i <= std_logic_vector(to_signed(integer( real(30)),WIDTH));
        midx_i <= std_logic_vector(to_signed(integer( real(42)),WIDTH));
        midy_i <= std_logic_vector(to_signed(integer( real(42)),WIDTH));
        
        --midx_i <= std_logic_vector(to_signed(integer( real(120)*real(2**FIXED_POINT_WIDTH)),WIDTH));
       -- midy_i <= std_logic_vector(to_signed(integer( real(120)*real(2**FIXED_POINT_WIDTH)),WIDTH));
       -- row_i <= std_logic_vector(to_signed(integer( real(54)*real(2**FIXED_POINT_WIDTH)),WIDTH));
       -- col_i <= std_logic_vector(to_signed(integer( real(22)*real(2**FIXED_POINT_WIDTH)),WIDTH));
        start_i <= '1';
       
        if ready_o /= '0' then
            wait until ready_o = '0';
        end if;
        wait for 200ns;
        start_i <= '0';
        if ready_o /= '1' then
            wait until ready_o = '1';
        end if;
        wait for 1000ns;
end process;
end Behavioral;
